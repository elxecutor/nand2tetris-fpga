/**
 * 1-bit register:
 * If load[t] == 1 then out[t+1] = in[t]
 *    else out does not change (out[t+1] = out[t])
 */

`default_nettype none
module Bit(
	input clk,
	input in,
	input load,
	output out
);

	// Put your code here:
	reg out_reg;
	always @(posedge clk) begin
		if (load) out_reg <= in;
	end
	assign out = out_reg;

endmodule
