/**
* 8-bit Shiftregister (shifts to left)
* if      (load == 1)  out[t+1] = in[t]
* else if (shift == 1) out[t+1] = out[t]<<1 | inLSB
* (shift one position to left and insert inLSB as least significant bit)
*/

`default_nettype none
module BitShift8L(
	input clk,
	input [7:0] in,
	input inLSB,
	input load,
	input shift,
	output [7:0] out
);

	// Put your code here:
	reg [7:0] out_reg;
	always @(posedge clk) begin
		if (load) out_reg <= in;
		else if (shift) out_reg <= {out_reg[6:0], inLSB};
		else out_reg <= out_reg;
	end
	assign out = out_reg;

endmodule
