/**
* RAM512 implements 512 Bytes of RAM addressed from 0 - 511
* out = M[address]
* if (load =i= 1) M[address][t+1] = in[t]
*/

`default_nettype none
module RAM512(
	input clk,
	input [8:0] address,
	input [15:0] in,
	input load,
	output [15:0] out
);
	
	// Put your code here:
	reg [15:0] mem [0:511];
	always @(posedge clk) begin
		if (load) mem[address] <= in;
	end
	assign out = mem[address];

endmodule
