/**
 * 16-bit register:
 * If load[t] == 1 then out[t+1] = in[t]
 * else out does not change
 */

`default_nettype none

module Register(
	input clk,
	input [15:0] in,
	input load,
	output [15:0] out
);

	// Put your code here:
	reg [15:0] out_reg;
	always @(posedge clk) begin
		if (load) out_reg <= in;
	end
	assign out = out_reg;

endmodule
